/* -------------------- REGMAP TEST -------------------------- */
$display("@ [TEST] Regmap Test started!");
/* ----------------------------------------------------------- */

    //| 1. Make a global reset;
    GlobalReset();

    //| Testing RW access for all RW registers