/* -------------------- RX/TX TEST -------------------------- */
$display("@ [TEST] RX/TX Test started!");
/* ----------------------------------------------------------- */

    //| 1. Make a global reset;
    GlobalReset();

    //| 2. Setup BAUDRATE and registers